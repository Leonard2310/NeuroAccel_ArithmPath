module datapath (A, B, opcode, Y, co);
  
  input signed [15:0] A, B;
  input [2:0] opcode;
  output signed [15:0] Y;
  output co;
  
  // add your code here
 
endmodule